// niosSys.v

// Generated using ACDS version 16.1 196

`timescale 1 ps / 1 ps
module niosSys (
		output wire [6:0]  hex_0_export,    //     hex_0.export
		output wire [6:0]  hex_1_export,    //     hex_1.export
		output wire [6:0]  hex_2_export,    //     hex_2.export
		output wire [6:0]  hex_3_export,    //     hex_3.export
		output wire [6:0]  hex_4_export,    //     hex_4.export
		output wire [6:0]  hex_5_export,    //     hex_5.export
		output wire [6:0]  hex_6_export,    //     hex_6.export
		output wire [6:0]  hex_7_export,    //     hex_7.export
		input  wire [3:0]  key_0_export,    //     key_0.export
		inout  wire [7:0]  lcd_DATA,        //       lcd.DATA
		output wire        lcd_ON,          //          .ON
		output wire        lcd_BLON,        //          .BLON
		output wire        lcd_EN,          //          .EN
		output wire        lcd_RS,          //          .RS
		output wire        lcd_RW,          //          .RW
		output wire [7:0]  ledg_export,     //      ledg.export
		output wire [17:0] leds_export,     //      leds.export
		input  wire        ref_clk_clk,     //   ref_clk.clk
		input  wire        ref_reset_reset, // ref_reset.reset
		inout  wire        sd_b_SD_cmd,     //        sd.b_SD_cmd
		inout  wire        sd_b_SD_dat,     //          .b_SD_dat
		inout  wire        sd_b_SD_dat3,    //          .b_SD_dat3
		output wire        sd_o_SD_clock,   //          .o_SD_clock
		output wire [12:0] sdram_addr,      //     sdram.addr
		output wire [1:0]  sdram_ba,        //          .ba
		output wire        sdram_cas_n,     //          .cas_n
		output wire        sdram_cke,       //          .cke
		output wire        sdram_cs_n,      //          .cs_n
		inout  wire [31:0] sdram_dq,        //          .dq
		output wire [3:0]  sdram_dqm,       //          .dqm
		output wire        sdram_ras_n,     //          .ras_n
		output wire        sdram_we_n,      //          .we_n
		output wire        sdram_clk_clk,   // sdram_clk.clk
		input  wire [17:0] switches_export  //  switches.export
	);

	wire         main_clk_sys_clk_clk;                                                                   // MAIN_CLK:sys_clk_clk -> [Altera_UP_SD_Card_Avalon_Interface_0:i_clock, HEX_0:clk, HEX_1:clk, HEX_2:clk, HEX_3:clk, HEX_4:clk, HEX_5:clk, HEX_6:clk, HEX_7:clk, High_Res_Timer:clk, KEY_0:clk, LEDG:clk, LEDs:clk, SDRAM:clk, Switches:clk, System_Clock_Timer:clk, TCM:clk, TCM:clk2, character_lcd_0:clk, irq_mapper:clk, jtag_uart_0:clk, mm_interconnect_0:MAIN_CLK_sys_clk_clk, mm_interconnect_1:MAIN_CLK_sys_clk_clk, myCPU:clk, rst_controller:clk, sysID:clock]
	wire  [31:0] mycpu_data_master_readdata;                                                             // mm_interconnect_0:myCPU_data_master_readdata -> myCPU:d_readdata
	wire         mycpu_data_master_waitrequest;                                                          // mm_interconnect_0:myCPU_data_master_waitrequest -> myCPU:d_waitrequest
	wire         mycpu_data_master_debugaccess;                                                          // myCPU:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:myCPU_data_master_debugaccess
	wire  [27:0] mycpu_data_master_address;                                                              // myCPU:d_address -> mm_interconnect_0:myCPU_data_master_address
	wire   [3:0] mycpu_data_master_byteenable;                                                           // myCPU:d_byteenable -> mm_interconnect_0:myCPU_data_master_byteenable
	wire         mycpu_data_master_read;                                                                 // myCPU:d_read -> mm_interconnect_0:myCPU_data_master_read
	wire         mycpu_data_master_readdatavalid;                                                        // mm_interconnect_0:myCPU_data_master_readdatavalid -> myCPU:d_readdatavalid
	wire         mycpu_data_master_write;                                                                // myCPU:d_write -> mm_interconnect_0:myCPU_data_master_write
	wire  [31:0] mycpu_data_master_writedata;                                                            // myCPU:d_writedata -> mm_interconnect_0:myCPU_data_master_writedata
	wire  [31:0] mycpu_instruction_master_readdata;                                                      // mm_interconnect_0:myCPU_instruction_master_readdata -> myCPU:i_readdata
	wire         mycpu_instruction_master_waitrequest;                                                   // mm_interconnect_0:myCPU_instruction_master_waitrequest -> myCPU:i_waitrequest
	wire  [27:0] mycpu_instruction_master_address;                                                       // myCPU:i_address -> mm_interconnect_0:myCPU_instruction_master_address
	wire         mycpu_instruction_master_read;                                                          // myCPU:i_read -> mm_interconnect_0:myCPU_instruction_master_read
	wire         mycpu_instruction_master_readdatavalid;                                                 // mm_interconnect_0:myCPU_instruction_master_readdatavalid -> myCPU:i_readdatavalid
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect;                             // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_chipselect -> jtag_uart_0:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata;                               // jtag_uart_0:av_readdata -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest;                            // jtag_uart_0:av_waitrequest -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address;                                // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_address -> jtag_uart_0:av_address
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read;                                   // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_read -> jtag_uart_0:av_read_n
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write;                                  // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_write -> jtag_uart_0:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata;                              // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_writedata -> jtag_uart_0:av_writedata
	wire         mm_interconnect_0_character_lcd_0_avalon_lcd_slave_chipselect;                          // mm_interconnect_0:character_lcd_0_avalon_lcd_slave_chipselect -> character_lcd_0:chipselect
	wire   [7:0] mm_interconnect_0_character_lcd_0_avalon_lcd_slave_readdata;                            // character_lcd_0:readdata -> mm_interconnect_0:character_lcd_0_avalon_lcd_slave_readdata
	wire         mm_interconnect_0_character_lcd_0_avalon_lcd_slave_waitrequest;                         // character_lcd_0:waitrequest -> mm_interconnect_0:character_lcd_0_avalon_lcd_slave_waitrequest
	wire   [0:0] mm_interconnect_0_character_lcd_0_avalon_lcd_slave_address;                             // mm_interconnect_0:character_lcd_0_avalon_lcd_slave_address -> character_lcd_0:address
	wire         mm_interconnect_0_character_lcd_0_avalon_lcd_slave_read;                                // mm_interconnect_0:character_lcd_0_avalon_lcd_slave_read -> character_lcd_0:read
	wire         mm_interconnect_0_character_lcd_0_avalon_lcd_slave_write;                               // mm_interconnect_0:character_lcd_0_avalon_lcd_slave_write -> character_lcd_0:write
	wire   [7:0] mm_interconnect_0_character_lcd_0_avalon_lcd_slave_writedata;                           // mm_interconnect_0:character_lcd_0_avalon_lcd_slave_writedata -> character_lcd_0:writedata
	wire         mm_interconnect_0_altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_chipselect;  // mm_interconnect_0:Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_chipselect -> Altera_UP_SD_Card_Avalon_Interface_0:i_avalon_chip_select
	wire  [31:0] mm_interconnect_0_altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_readdata;    // Altera_UP_SD_Card_Avalon_Interface_0:o_avalon_readdata -> mm_interconnect_0:Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_readdata
	wire         mm_interconnect_0_altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_waitrequest; // Altera_UP_SD_Card_Avalon_Interface_0:o_avalon_waitrequest -> mm_interconnect_0:Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_waitrequest
	wire   [7:0] mm_interconnect_0_altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_address;     // mm_interconnect_0:Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_address -> Altera_UP_SD_Card_Avalon_Interface_0:i_avalon_address
	wire         mm_interconnect_0_altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_read;        // mm_interconnect_0:Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_read -> Altera_UP_SD_Card_Avalon_Interface_0:i_avalon_read
	wire   [3:0] mm_interconnect_0_altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_byteenable;  // mm_interconnect_0:Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_byteenable -> Altera_UP_SD_Card_Avalon_Interface_0:i_avalon_byteenable
	wire         mm_interconnect_0_altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_write;       // mm_interconnect_0:Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_write -> Altera_UP_SD_Card_Avalon_Interface_0:i_avalon_write
	wire  [31:0] mm_interconnect_0_altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_writedata;   // mm_interconnect_0:Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_writedata -> Altera_UP_SD_Card_Avalon_Interface_0:i_avalon_writedata
	wire  [31:0] mm_interconnect_0_sysid_control_slave_readdata;                                         // sysID:readdata -> mm_interconnect_0:sysID_control_slave_readdata
	wire   [0:0] mm_interconnect_0_sysid_control_slave_address;                                          // mm_interconnect_0:sysID_control_slave_address -> sysID:address
	wire  [31:0] mm_interconnect_0_mycpu_debug_mem_slave_readdata;                                       // myCPU:debug_mem_slave_readdata -> mm_interconnect_0:myCPU_debug_mem_slave_readdata
	wire         mm_interconnect_0_mycpu_debug_mem_slave_waitrequest;                                    // myCPU:debug_mem_slave_waitrequest -> mm_interconnect_0:myCPU_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_mycpu_debug_mem_slave_debugaccess;                                    // mm_interconnect_0:myCPU_debug_mem_slave_debugaccess -> myCPU:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_mycpu_debug_mem_slave_address;                                        // mm_interconnect_0:myCPU_debug_mem_slave_address -> myCPU:debug_mem_slave_address
	wire         mm_interconnect_0_mycpu_debug_mem_slave_read;                                           // mm_interconnect_0:myCPU_debug_mem_slave_read -> myCPU:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_mycpu_debug_mem_slave_byteenable;                                     // mm_interconnect_0:myCPU_debug_mem_slave_byteenable -> myCPU:debug_mem_slave_byteenable
	wire         mm_interconnect_0_mycpu_debug_mem_slave_write;                                          // mm_interconnect_0:myCPU_debug_mem_slave_write -> myCPU:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_mycpu_debug_mem_slave_writedata;                                      // mm_interconnect_0:myCPU_debug_mem_slave_writedata -> myCPU:debug_mem_slave_writedata
	wire         mm_interconnect_0_system_clock_timer_s1_chipselect;                                     // mm_interconnect_0:System_Clock_Timer_s1_chipselect -> System_Clock_Timer:chipselect
	wire  [15:0] mm_interconnect_0_system_clock_timer_s1_readdata;                                       // System_Clock_Timer:readdata -> mm_interconnect_0:System_Clock_Timer_s1_readdata
	wire   [2:0] mm_interconnect_0_system_clock_timer_s1_address;                                        // mm_interconnect_0:System_Clock_Timer_s1_address -> System_Clock_Timer:address
	wire         mm_interconnect_0_system_clock_timer_s1_write;                                          // mm_interconnect_0:System_Clock_Timer_s1_write -> System_Clock_Timer:write_n
	wire  [15:0] mm_interconnect_0_system_clock_timer_s1_writedata;                                      // mm_interconnect_0:System_Clock_Timer_s1_writedata -> System_Clock_Timer:writedata
	wire         mm_interconnect_0_high_res_timer_s1_chipselect;                                         // mm_interconnect_0:High_Res_Timer_s1_chipselect -> High_Res_Timer:chipselect
	wire  [15:0] mm_interconnect_0_high_res_timer_s1_readdata;                                           // High_Res_Timer:readdata -> mm_interconnect_0:High_Res_Timer_s1_readdata
	wire   [2:0] mm_interconnect_0_high_res_timer_s1_address;                                            // mm_interconnect_0:High_Res_Timer_s1_address -> High_Res_Timer:address
	wire         mm_interconnect_0_high_res_timer_s1_write;                                              // mm_interconnect_0:High_Res_Timer_s1_write -> High_Res_Timer:write_n
	wire  [15:0] mm_interconnect_0_high_res_timer_s1_writedata;                                          // mm_interconnect_0:High_Res_Timer_s1_writedata -> High_Res_Timer:writedata
	wire         mm_interconnect_0_switches_s1_chipselect;                                               // mm_interconnect_0:Switches_s1_chipselect -> Switches:chipselect
	wire  [31:0] mm_interconnect_0_switches_s1_readdata;                                                 // Switches:readdata -> mm_interconnect_0:Switches_s1_readdata
	wire   [1:0] mm_interconnect_0_switches_s1_address;                                                  // mm_interconnect_0:Switches_s1_address -> Switches:address
	wire         mm_interconnect_0_switches_s1_write;                                                    // mm_interconnect_0:Switches_s1_write -> Switches:write_n
	wire  [31:0] mm_interconnect_0_switches_s1_writedata;                                                // mm_interconnect_0:Switches_s1_writedata -> Switches:writedata
	wire         mm_interconnect_0_leds_s1_chipselect;                                                   // mm_interconnect_0:LEDs_s1_chipselect -> LEDs:chipselect
	wire  [31:0] mm_interconnect_0_leds_s1_readdata;                                                     // LEDs:readdata -> mm_interconnect_0:LEDs_s1_readdata
	wire   [1:0] mm_interconnect_0_leds_s1_address;                                                      // mm_interconnect_0:LEDs_s1_address -> LEDs:address
	wire         mm_interconnect_0_leds_s1_write;                                                        // mm_interconnect_0:LEDs_s1_write -> LEDs:write_n
	wire  [31:0] mm_interconnect_0_leds_s1_writedata;                                                    // mm_interconnect_0:LEDs_s1_writedata -> LEDs:writedata
	wire         mm_interconnect_0_hex_0_s1_chipselect;                                                  // mm_interconnect_0:HEX_0_s1_chipselect -> HEX_0:chipselect
	wire  [31:0] mm_interconnect_0_hex_0_s1_readdata;                                                    // HEX_0:readdata -> mm_interconnect_0:HEX_0_s1_readdata
	wire   [1:0] mm_interconnect_0_hex_0_s1_address;                                                     // mm_interconnect_0:HEX_0_s1_address -> HEX_0:address
	wire         mm_interconnect_0_hex_0_s1_write;                                                       // mm_interconnect_0:HEX_0_s1_write -> HEX_0:write_n
	wire  [31:0] mm_interconnect_0_hex_0_s1_writedata;                                                   // mm_interconnect_0:HEX_0_s1_writedata -> HEX_0:writedata
	wire         mm_interconnect_0_hex_1_s1_chipselect;                                                  // mm_interconnect_0:HEX_1_s1_chipselect -> HEX_1:chipselect
	wire  [31:0] mm_interconnect_0_hex_1_s1_readdata;                                                    // HEX_1:readdata -> mm_interconnect_0:HEX_1_s1_readdata
	wire   [1:0] mm_interconnect_0_hex_1_s1_address;                                                     // mm_interconnect_0:HEX_1_s1_address -> HEX_1:address
	wire         mm_interconnect_0_hex_1_s1_write;                                                       // mm_interconnect_0:HEX_1_s1_write -> HEX_1:write_n
	wire  [31:0] mm_interconnect_0_hex_1_s1_writedata;                                                   // mm_interconnect_0:HEX_1_s1_writedata -> HEX_1:writedata
	wire         mm_interconnect_0_hex_2_s1_chipselect;                                                  // mm_interconnect_0:HEX_2_s1_chipselect -> HEX_2:chipselect
	wire  [31:0] mm_interconnect_0_hex_2_s1_readdata;                                                    // HEX_2:readdata -> mm_interconnect_0:HEX_2_s1_readdata
	wire   [1:0] mm_interconnect_0_hex_2_s1_address;                                                     // mm_interconnect_0:HEX_2_s1_address -> HEX_2:address
	wire         mm_interconnect_0_hex_2_s1_write;                                                       // mm_interconnect_0:HEX_2_s1_write -> HEX_2:write_n
	wire  [31:0] mm_interconnect_0_hex_2_s1_writedata;                                                   // mm_interconnect_0:HEX_2_s1_writedata -> HEX_2:writedata
	wire         mm_interconnect_0_hex_3_s1_chipselect;                                                  // mm_interconnect_0:HEX_3_s1_chipselect -> HEX_3:chipselect
	wire  [31:0] mm_interconnect_0_hex_3_s1_readdata;                                                    // HEX_3:readdata -> mm_interconnect_0:HEX_3_s1_readdata
	wire   [1:0] mm_interconnect_0_hex_3_s1_address;                                                     // mm_interconnect_0:HEX_3_s1_address -> HEX_3:address
	wire         mm_interconnect_0_hex_3_s1_write;                                                       // mm_interconnect_0:HEX_3_s1_write -> HEX_3:write_n
	wire  [31:0] mm_interconnect_0_hex_3_s1_writedata;                                                   // mm_interconnect_0:HEX_3_s1_writedata -> HEX_3:writedata
	wire         mm_interconnect_0_hex_4_s1_chipselect;                                                  // mm_interconnect_0:HEX_4_s1_chipselect -> HEX_4:chipselect
	wire  [31:0] mm_interconnect_0_hex_4_s1_readdata;                                                    // HEX_4:readdata -> mm_interconnect_0:HEX_4_s1_readdata
	wire   [1:0] mm_interconnect_0_hex_4_s1_address;                                                     // mm_interconnect_0:HEX_4_s1_address -> HEX_4:address
	wire         mm_interconnect_0_hex_4_s1_write;                                                       // mm_interconnect_0:HEX_4_s1_write -> HEX_4:write_n
	wire  [31:0] mm_interconnect_0_hex_4_s1_writedata;                                                   // mm_interconnect_0:HEX_4_s1_writedata -> HEX_4:writedata
	wire         mm_interconnect_0_hex_5_s1_chipselect;                                                  // mm_interconnect_0:HEX_5_s1_chipselect -> HEX_5:chipselect
	wire  [31:0] mm_interconnect_0_hex_5_s1_readdata;                                                    // HEX_5:readdata -> mm_interconnect_0:HEX_5_s1_readdata
	wire   [1:0] mm_interconnect_0_hex_5_s1_address;                                                     // mm_interconnect_0:HEX_5_s1_address -> HEX_5:address
	wire         mm_interconnect_0_hex_5_s1_write;                                                       // mm_interconnect_0:HEX_5_s1_write -> HEX_5:write_n
	wire  [31:0] mm_interconnect_0_hex_5_s1_writedata;                                                   // mm_interconnect_0:HEX_5_s1_writedata -> HEX_5:writedata
	wire         mm_interconnect_0_hex_6_s1_chipselect;                                                  // mm_interconnect_0:HEX_6_s1_chipselect -> HEX_6:chipselect
	wire  [31:0] mm_interconnect_0_hex_6_s1_readdata;                                                    // HEX_6:readdata -> mm_interconnect_0:HEX_6_s1_readdata
	wire   [1:0] mm_interconnect_0_hex_6_s1_address;                                                     // mm_interconnect_0:HEX_6_s1_address -> HEX_6:address
	wire         mm_interconnect_0_hex_6_s1_write;                                                       // mm_interconnect_0:HEX_6_s1_write -> HEX_6:write_n
	wire  [31:0] mm_interconnect_0_hex_6_s1_writedata;                                                   // mm_interconnect_0:HEX_6_s1_writedata -> HEX_6:writedata
	wire         mm_interconnect_0_hex_7_s1_chipselect;                                                  // mm_interconnect_0:HEX_7_s1_chipselect -> HEX_7:chipselect
	wire  [31:0] mm_interconnect_0_hex_7_s1_readdata;                                                    // HEX_7:readdata -> mm_interconnect_0:HEX_7_s1_readdata
	wire   [1:0] mm_interconnect_0_hex_7_s1_address;                                                     // mm_interconnect_0:HEX_7_s1_address -> HEX_7:address
	wire         mm_interconnect_0_hex_7_s1_write;                                                       // mm_interconnect_0:HEX_7_s1_write -> HEX_7:write_n
	wire  [31:0] mm_interconnect_0_hex_7_s1_writedata;                                                   // mm_interconnect_0:HEX_7_s1_writedata -> HEX_7:writedata
	wire         mm_interconnect_0_ledg_s1_chipselect;                                                   // mm_interconnect_0:LEDG_s1_chipselect -> LEDG:chipselect
	wire  [31:0] mm_interconnect_0_ledg_s1_readdata;                                                     // LEDG:readdata -> mm_interconnect_0:LEDG_s1_readdata
	wire   [1:0] mm_interconnect_0_ledg_s1_address;                                                      // mm_interconnect_0:LEDG_s1_address -> LEDG:address
	wire         mm_interconnect_0_ledg_s1_write;                                                        // mm_interconnect_0:LEDG_s1_write -> LEDG:write_n
	wire  [31:0] mm_interconnect_0_ledg_s1_writedata;                                                    // mm_interconnect_0:LEDG_s1_writedata -> LEDG:writedata
	wire         mm_interconnect_0_key_0_s1_chipselect;                                                  // mm_interconnect_0:KEY_0_s1_chipselect -> KEY_0:chipselect
	wire  [31:0] mm_interconnect_0_key_0_s1_readdata;                                                    // KEY_0:readdata -> mm_interconnect_0:KEY_0_s1_readdata
	wire   [1:0] mm_interconnect_0_key_0_s1_address;                                                     // mm_interconnect_0:KEY_0_s1_address -> KEY_0:address
	wire         mm_interconnect_0_key_0_s1_write;                                                       // mm_interconnect_0:KEY_0_s1_write -> KEY_0:write_n
	wire  [31:0] mm_interconnect_0_key_0_s1_writedata;                                                   // mm_interconnect_0:KEY_0_s1_writedata -> KEY_0:writedata
	wire         mm_interconnect_0_sdram_s1_chipselect;                                                  // mm_interconnect_0:SDRAM_s1_chipselect -> SDRAM:az_cs
	wire  [31:0] mm_interconnect_0_sdram_s1_readdata;                                                    // SDRAM:za_data -> mm_interconnect_0:SDRAM_s1_readdata
	wire         mm_interconnect_0_sdram_s1_waitrequest;                                                 // SDRAM:za_waitrequest -> mm_interconnect_0:SDRAM_s1_waitrequest
	wire  [24:0] mm_interconnect_0_sdram_s1_address;                                                     // mm_interconnect_0:SDRAM_s1_address -> SDRAM:az_addr
	wire         mm_interconnect_0_sdram_s1_read;                                                        // mm_interconnect_0:SDRAM_s1_read -> SDRAM:az_rd_n
	wire   [3:0] mm_interconnect_0_sdram_s1_byteenable;                                                  // mm_interconnect_0:SDRAM_s1_byteenable -> SDRAM:az_be_n
	wire         mm_interconnect_0_sdram_s1_readdatavalid;                                               // SDRAM:za_valid -> mm_interconnect_0:SDRAM_s1_readdatavalid
	wire         mm_interconnect_0_sdram_s1_write;                                                       // mm_interconnect_0:SDRAM_s1_write -> SDRAM:az_wr_n
	wire  [31:0] mm_interconnect_0_sdram_s1_writedata;                                                   // mm_interconnect_0:SDRAM_s1_writedata -> SDRAM:az_data
	wire         mm_interconnect_0_tcm_s2_chipselect;                                                    // mm_interconnect_0:TCM_s2_chipselect -> TCM:chipselect2
	wire  [31:0] mm_interconnect_0_tcm_s2_readdata;                                                      // TCM:readdata2 -> mm_interconnect_0:TCM_s2_readdata
	wire   [8:0] mm_interconnect_0_tcm_s2_address;                                                       // mm_interconnect_0:TCM_s2_address -> TCM:address2
	wire   [3:0] mm_interconnect_0_tcm_s2_byteenable;                                                    // mm_interconnect_0:TCM_s2_byteenable -> TCM:byteenable2
	wire         mm_interconnect_0_tcm_s2_write;                                                         // mm_interconnect_0:TCM_s2_write -> TCM:write2
	wire  [31:0] mm_interconnect_0_tcm_s2_writedata;                                                     // mm_interconnect_0:TCM_s2_writedata -> TCM:writedata2
	wire         mm_interconnect_0_tcm_s2_clken;                                                         // mm_interconnect_0:TCM_s2_clken -> TCM:clken2
	wire  [31:0] mycpu_tightly_coupled_instruction_master_0_readdata;                                    // mm_interconnect_1:myCPU_tightly_coupled_instruction_master_0_readdata -> myCPU:itcm0_readdata
	wire  [10:0] mycpu_tightly_coupled_instruction_master_0_address;                                     // myCPU:itcm0_address -> mm_interconnect_1:myCPU_tightly_coupled_instruction_master_0_address
	wire         mycpu_tightly_coupled_instruction_master_0_read;                                        // myCPU:itcm0_read -> mm_interconnect_1:myCPU_tightly_coupled_instruction_master_0_read
	wire         mycpu_tightly_coupled_instruction_master_0_clken;                                       // myCPU:itcm0_clken -> mm_interconnect_1:myCPU_tightly_coupled_instruction_master_0_clken
	wire         mm_interconnect_1_tcm_s1_chipselect;                                                    // mm_interconnect_1:TCM_s1_chipselect -> TCM:chipselect
	wire  [31:0] mm_interconnect_1_tcm_s1_readdata;                                                      // TCM:readdata -> mm_interconnect_1:TCM_s1_readdata
	wire   [8:0] mm_interconnect_1_tcm_s1_address;                                                       // mm_interconnect_1:TCM_s1_address -> TCM:address
	wire   [3:0] mm_interconnect_1_tcm_s1_byteenable;                                                    // mm_interconnect_1:TCM_s1_byteenable -> TCM:byteenable
	wire         mm_interconnect_1_tcm_s1_write;                                                         // mm_interconnect_1:TCM_s1_write -> TCM:write
	wire  [31:0] mm_interconnect_1_tcm_s1_writedata;                                                     // mm_interconnect_1:TCM_s1_writedata -> TCM:writedata
	wire         mm_interconnect_1_tcm_s1_clken;                                                         // mm_interconnect_1:TCM_s1_clken -> TCM:clken
	wire         irq_mapper_receiver0_irq;                                                               // jtag_uart_0:av_irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                                               // System_Clock_Timer:irq -> irq_mapper:receiver1_irq
	wire         irq_mapper_receiver2_irq;                                                               // High_Res_Timer:irq -> irq_mapper:receiver2_irq
	wire         irq_mapper_receiver3_irq;                                                               // Switches:irq -> irq_mapper:receiver3_irq
	wire         irq_mapper_receiver4_irq;                                                               // KEY_0:irq -> irq_mapper:receiver4_irq
	wire  [31:0] mycpu_irq_irq;                                                                          // irq_mapper:sender_irq -> myCPU:irq
	wire         rst_controller_reset_out_reset;                                                         // rst_controller:reset_out -> [Altera_UP_SD_Card_Avalon_Interface_0:i_reset_n, HEX_0:reset_n, HEX_1:reset_n, HEX_2:reset_n, HEX_3:reset_n, HEX_4:reset_n, HEX_5:reset_n, HEX_6:reset_n, HEX_7:reset_n, High_Res_Timer:reset_n, KEY_0:reset_n, LEDG:reset_n, LEDs:reset_n, SDRAM:reset_n, Switches:reset_n, System_Clock_Timer:reset_n, TCM:reset, TCM:reset2, character_lcd_0:reset, irq_mapper:reset, jtag_uart_0:rst_n, mm_interconnect_0:myCPU_reset_reset_bridge_in_reset_reset, mm_interconnect_1:myCPU_reset_reset_bridge_in_reset_reset, myCPU:reset_n, rst_translator:in_reset, sysID:reset_n]
	wire         rst_controller_reset_out_reset_req;                                                     // rst_controller:reset_req -> [TCM:reset_req, TCM:reset_req2, myCPU:reset_req, rst_translator:reset_req_in]
	wire         mycpu_debug_reset_request_reset;                                                        // myCPU:debug_reset_request -> rst_controller:reset_in0
	wire         main_clk_reset_source_reset;                                                            // MAIN_CLK:reset_source_reset -> rst_controller:reset_in1

	Altera_UP_SD_Card_Avalon_Interface altera_up_sd_card_avalon_interface_0 (
		.i_avalon_chip_select (mm_interconnect_0_altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_chipselect),  // avalon_sdcard_slave.chipselect
		.i_avalon_address     (mm_interconnect_0_altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_address),     //                    .address
		.i_avalon_read        (mm_interconnect_0_altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_read),        //                    .read
		.i_avalon_write       (mm_interconnect_0_altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_write),       //                    .write
		.i_avalon_byteenable  (mm_interconnect_0_altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_byteenable),  //                    .byteenable
		.i_avalon_writedata   (mm_interconnect_0_altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_writedata),   //                    .writedata
		.o_avalon_readdata    (mm_interconnect_0_altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_readdata),    //                    .readdata
		.o_avalon_waitrequest (mm_interconnect_0_altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_waitrequest), //                    .waitrequest
		.i_clock              (main_clk_sys_clk_clk),                                                                   //                 clk.clk
		.i_reset_n            (~rst_controller_reset_out_reset),                                                        //               reset.reset_n
		.b_SD_cmd             (sd_b_SD_cmd),                                                                            //         conduit_end.export
		.b_SD_dat             (sd_b_SD_dat),                                                                            //                    .export
		.b_SD_dat3            (sd_b_SD_dat3),                                                                           //                    .export
		.o_SD_clock           (sd_o_SD_clock)                                                                           //                    .export
	);

	niosSys_HEX_0 hex_0 (
		.clk        (main_clk_sys_clk_clk),                  //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_hex_0_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_hex_0_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_hex_0_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_hex_0_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_hex_0_s1_readdata),   //                    .readdata
		.out_port   (hex_0_export)                           // external_connection.export
	);

	niosSys_HEX_0 hex_1 (
		.clk        (main_clk_sys_clk_clk),                  //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_hex_1_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_hex_1_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_hex_1_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_hex_1_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_hex_1_s1_readdata),   //                    .readdata
		.out_port   (hex_1_export)                           // external_connection.export
	);

	niosSys_HEX_0 hex_2 (
		.clk        (main_clk_sys_clk_clk),                  //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_hex_2_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_hex_2_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_hex_2_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_hex_2_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_hex_2_s1_readdata),   //                    .readdata
		.out_port   (hex_2_export)                           // external_connection.export
	);

	niosSys_HEX_0 hex_3 (
		.clk        (main_clk_sys_clk_clk),                  //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_hex_3_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_hex_3_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_hex_3_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_hex_3_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_hex_3_s1_readdata),   //                    .readdata
		.out_port   (hex_3_export)                           // external_connection.export
	);

	niosSys_HEX_0 hex_4 (
		.clk        (main_clk_sys_clk_clk),                  //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_hex_4_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_hex_4_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_hex_4_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_hex_4_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_hex_4_s1_readdata),   //                    .readdata
		.out_port   (hex_4_export)                           // external_connection.export
	);

	niosSys_HEX_0 hex_5 (
		.clk        (main_clk_sys_clk_clk),                  //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_hex_5_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_hex_5_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_hex_5_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_hex_5_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_hex_5_s1_readdata),   //                    .readdata
		.out_port   (hex_5_export)                           // external_connection.export
	);

	niosSys_HEX_0 hex_6 (
		.clk        (main_clk_sys_clk_clk),                  //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_hex_6_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_hex_6_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_hex_6_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_hex_6_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_hex_6_s1_readdata),   //                    .readdata
		.out_port   (hex_6_export)                           // external_connection.export
	);

	niosSys_HEX_0 hex_7 (
		.clk        (main_clk_sys_clk_clk),                  //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_hex_7_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_hex_7_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_hex_7_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_hex_7_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_hex_7_s1_readdata),   //                    .readdata
		.out_port   (hex_7_export)                           // external_connection.export
	);

	niosSys_High_Res_Timer high_res_timer (
		.clk        (main_clk_sys_clk_clk),                           //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                // reset.reset_n
		.address    (mm_interconnect_0_high_res_timer_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_high_res_timer_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_high_res_timer_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_high_res_timer_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_high_res_timer_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver2_irq)                        //   irq.irq
	);

	niosSys_KEY_0 key_0 (
		.clk        (main_clk_sys_clk_clk),                  //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_key_0_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_key_0_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_key_0_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_key_0_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_key_0_s1_readdata),   //                    .readdata
		.in_port    (key_0_export),                          // external_connection.export
		.irq        (irq_mapper_receiver4_irq)               //                 irq.irq
	);

	niosSys_LEDG ledg (
		.clk        (main_clk_sys_clk_clk),                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_ledg_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_ledg_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_ledg_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_ledg_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_ledg_s1_readdata),   //                    .readdata
		.out_port   (ledg_export)                           // external_connection.export
	);

	niosSys_LEDs leds (
		.clk        (main_clk_sys_clk_clk),                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_leds_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_leds_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_leds_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_leds_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_leds_s1_readdata),   //                    .readdata
		.out_port   (leds_export)                           // external_connection.export
	);

	niosSys_MAIN_CLK main_clk (
		.ref_clk_clk        (ref_clk_clk),                 //      ref_clk.clk
		.ref_reset_reset    (ref_reset_reset),             //    ref_reset.reset
		.sys_clk_clk        (main_clk_sys_clk_clk),        //      sys_clk.clk
		.sdram_clk_clk      (sdram_clk_clk),               //    sdram_clk.clk
		.reset_source_reset (main_clk_reset_source_reset)  // reset_source.reset
	);

	niosSys_SDRAM sdram (
		.clk            (main_clk_sys_clk_clk),                     //   clk.clk
		.reset_n        (~rst_controller_reset_out_reset),          // reset.reset_n
		.az_addr        (mm_interconnect_0_sdram_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_0_sdram_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_0_sdram_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_0_sdram_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_0_sdram_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_0_sdram_s1_write),        //      .write_n
		.za_data        (mm_interconnect_0_sdram_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_0_sdram_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_0_sdram_s1_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_addr),                               //  wire.export
		.zs_ba          (sdram_ba),                                 //      .export
		.zs_cas_n       (sdram_cas_n),                              //      .export
		.zs_cke         (sdram_cke),                                //      .export
		.zs_cs_n        (sdram_cs_n),                               //      .export
		.zs_dq          (sdram_dq),                                 //      .export
		.zs_dqm         (sdram_dqm),                                //      .export
		.zs_ras_n       (sdram_ras_n),                              //      .export
		.zs_we_n        (sdram_we_n)                                //      .export
	);

	niosSys_Switches switches (
		.clk        (main_clk_sys_clk_clk),                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address    (mm_interconnect_0_switches_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_switches_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_switches_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_switches_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_switches_s1_readdata),   //                    .readdata
		.in_port    (switches_export),                          // external_connection.export
		.irq        (irq_mapper_receiver3_irq)                  //                 irq.irq
	);

	niosSys_High_Res_Timer system_clock_timer (
		.clk        (main_clk_sys_clk_clk),                               //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                    // reset.reset_n
		.address    (mm_interconnect_0_system_clock_timer_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_system_clock_timer_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_system_clock_timer_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_system_clock_timer_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_system_clock_timer_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver1_irq)                            //   irq.irq
	);

	niosSys_TCM tcm (
		.clk         (main_clk_sys_clk_clk),                //   clk1.clk
		.address     (mm_interconnect_1_tcm_s1_address),    //     s1.address
		.clken       (mm_interconnect_1_tcm_s1_clken),      //       .clken
		.chipselect  (mm_interconnect_1_tcm_s1_chipselect), //       .chipselect
		.write       (mm_interconnect_1_tcm_s1_write),      //       .write
		.readdata    (mm_interconnect_1_tcm_s1_readdata),   //       .readdata
		.writedata   (mm_interconnect_1_tcm_s1_writedata),  //       .writedata
		.byteenable  (mm_interconnect_1_tcm_s1_byteenable), //       .byteenable
		.reset       (rst_controller_reset_out_reset),      // reset1.reset
		.reset_req   (rst_controller_reset_out_reset_req),  //       .reset_req
		.address2    (mm_interconnect_0_tcm_s2_address),    //     s2.address
		.chipselect2 (mm_interconnect_0_tcm_s2_chipselect), //       .chipselect
		.clken2      (mm_interconnect_0_tcm_s2_clken),      //       .clken
		.write2      (mm_interconnect_0_tcm_s2_write),      //       .write
		.readdata2   (mm_interconnect_0_tcm_s2_readdata),   //       .readdata
		.writedata2  (mm_interconnect_0_tcm_s2_writedata),  //       .writedata
		.byteenable2 (mm_interconnect_0_tcm_s2_byteenable), //       .byteenable
		.clk2        (main_clk_sys_clk_clk),                //   clk2.clk
		.reset2      (rst_controller_reset_out_reset),      // reset2.reset
		.reset_req2  (rst_controller_reset_out_reset_req),  //       .reset_req
		.freeze      (1'b0)                                 // (terminated)
	);

	niosSys_character_lcd_0 character_lcd_0 (
		.clk         (main_clk_sys_clk_clk),                                           //                clk.clk
		.reset       (rst_controller_reset_out_reset),                                 //              reset.reset
		.address     (mm_interconnect_0_character_lcd_0_avalon_lcd_slave_address),     //   avalon_lcd_slave.address
		.chipselect  (mm_interconnect_0_character_lcd_0_avalon_lcd_slave_chipselect),  //                   .chipselect
		.read        (mm_interconnect_0_character_lcd_0_avalon_lcd_slave_read),        //                   .read
		.write       (mm_interconnect_0_character_lcd_0_avalon_lcd_slave_write),       //                   .write
		.writedata   (mm_interconnect_0_character_lcd_0_avalon_lcd_slave_writedata),   //                   .writedata
		.readdata    (mm_interconnect_0_character_lcd_0_avalon_lcd_slave_readdata),    //                   .readdata
		.waitrequest (mm_interconnect_0_character_lcd_0_avalon_lcd_slave_waitrequest), //                   .waitrequest
		.LCD_DATA    (lcd_DATA),                                                       // external_interface.export
		.LCD_ON      (lcd_ON),                                                         //                   .export
		.LCD_BLON    (lcd_BLON),                                                       //                   .export
		.LCD_EN      (lcd_EN),                                                         //                   .export
		.LCD_RS      (lcd_RS),                                                         //                   .export
		.LCD_RW      (lcd_RW)                                                          //                   .export
	);

	niosSys_jtag_uart_0 jtag_uart_0 (
		.clk            (main_clk_sys_clk_clk),                                        //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                             //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                     //               irq.irq
	);

	niosSys_myCPU mycpu (
		.clk                                 (main_clk_sys_clk_clk),                                //                                  clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                     //                                reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                  //                                     .reset_req
		.d_address                           (mycpu_data_master_address),                           //                          data_master.address
		.d_byteenable                        (mycpu_data_master_byteenable),                        //                                     .byteenable
		.d_read                              (mycpu_data_master_read),                              //                                     .read
		.d_readdata                          (mycpu_data_master_readdata),                          //                                     .readdata
		.d_waitrequest                       (mycpu_data_master_waitrequest),                       //                                     .waitrequest
		.d_write                             (mycpu_data_master_write),                             //                                     .write
		.d_writedata                         (mycpu_data_master_writedata),                         //                                     .writedata
		.d_readdatavalid                     (mycpu_data_master_readdatavalid),                     //                                     .readdatavalid
		.debug_mem_slave_debugaccess_to_roms (mycpu_data_master_debugaccess),                       //                                     .debugaccess
		.i_address                           (mycpu_instruction_master_address),                    //                   instruction_master.address
		.i_read                              (mycpu_instruction_master_read),                       //                                     .read
		.i_readdata                          (mycpu_instruction_master_readdata),                   //                                     .readdata
		.i_waitrequest                       (mycpu_instruction_master_waitrequest),                //                                     .waitrequest
		.i_readdatavalid                     (mycpu_instruction_master_readdatavalid),              //                                     .readdatavalid
		.itcm0_readdata                      (mycpu_tightly_coupled_instruction_master_0_readdata), // tightly_coupled_instruction_master_0.readdata
		.itcm0_address                       (mycpu_tightly_coupled_instruction_master_0_address),  //                                     .address
		.itcm0_read                          (mycpu_tightly_coupled_instruction_master_0_read),     //                                     .read
		.itcm0_clken                         (mycpu_tightly_coupled_instruction_master_0_clken),    //                                     .clken
		.irq                                 (mycpu_irq_irq),                                       //                                  irq.irq
		.debug_reset_request                 (mycpu_debug_reset_request_reset),                     //                  debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_mycpu_debug_mem_slave_address),     //                      debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_mycpu_debug_mem_slave_byteenable),  //                                     .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_mycpu_debug_mem_slave_debugaccess), //                                     .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_mycpu_debug_mem_slave_read),        //                                     .read
		.debug_mem_slave_readdata            (mm_interconnect_0_mycpu_debug_mem_slave_readdata),    //                                     .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_mycpu_debug_mem_slave_waitrequest), //                                     .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_mycpu_debug_mem_slave_write),       //                                     .write
		.debug_mem_slave_writedata           (mm_interconnect_0_mycpu_debug_mem_slave_writedata),   //                                     .writedata
		.dummy_ci_port                       ()                                                     //            custom_instruction_master.readra
	);

	niosSys_sysID sysid (
		.clock    (main_clk_sys_clk_clk),                           //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_control_slave_address)   //              .address
	);

	niosSys_mm_interconnect_0 mm_interconnect_0 (
		.MAIN_CLK_sys_clk_clk                                                 (main_clk_sys_clk_clk),                                                                   //                                         MAIN_CLK_sys_clk.clk
		.myCPU_reset_reset_bridge_in_reset_reset                              (rst_controller_reset_out_reset),                                                         //                        myCPU_reset_reset_bridge_in_reset.reset
		.myCPU_data_master_address                                            (mycpu_data_master_address),                                                              //                                        myCPU_data_master.address
		.myCPU_data_master_waitrequest                                        (mycpu_data_master_waitrequest),                                                          //                                                         .waitrequest
		.myCPU_data_master_byteenable                                         (mycpu_data_master_byteenable),                                                           //                                                         .byteenable
		.myCPU_data_master_read                                               (mycpu_data_master_read),                                                                 //                                                         .read
		.myCPU_data_master_readdata                                           (mycpu_data_master_readdata),                                                             //                                                         .readdata
		.myCPU_data_master_readdatavalid                                      (mycpu_data_master_readdatavalid),                                                        //                                                         .readdatavalid
		.myCPU_data_master_write                                              (mycpu_data_master_write),                                                                //                                                         .write
		.myCPU_data_master_writedata                                          (mycpu_data_master_writedata),                                                            //                                                         .writedata
		.myCPU_data_master_debugaccess                                        (mycpu_data_master_debugaccess),                                                          //                                                         .debugaccess
		.myCPU_instruction_master_address                                     (mycpu_instruction_master_address),                                                       //                                 myCPU_instruction_master.address
		.myCPU_instruction_master_waitrequest                                 (mycpu_instruction_master_waitrequest),                                                   //                                                         .waitrequest
		.myCPU_instruction_master_read                                        (mycpu_instruction_master_read),                                                          //                                                         .read
		.myCPU_instruction_master_readdata                                    (mycpu_instruction_master_readdata),                                                      //                                                         .readdata
		.myCPU_instruction_master_readdatavalid                               (mycpu_instruction_master_readdatavalid),                                                 //                                                         .readdatavalid
		.Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_address     (mm_interconnect_0_altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_address),     // Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave.address
		.Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_write       (mm_interconnect_0_altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_write),       //                                                         .write
		.Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_read        (mm_interconnect_0_altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_read),        //                                                         .read
		.Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_readdata    (mm_interconnect_0_altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_readdata),    //                                                         .readdata
		.Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_writedata   (mm_interconnect_0_altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_writedata),   //                                                         .writedata
		.Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_byteenable  (mm_interconnect_0_altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_byteenable),  //                                                         .byteenable
		.Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_waitrequest (mm_interconnect_0_altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_waitrequest), //                                                         .waitrequest
		.Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_chipselect  (mm_interconnect_0_altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_chipselect),  //                                                         .chipselect
		.character_lcd_0_avalon_lcd_slave_address                             (mm_interconnect_0_character_lcd_0_avalon_lcd_slave_address),                             //                         character_lcd_0_avalon_lcd_slave.address
		.character_lcd_0_avalon_lcd_slave_write                               (mm_interconnect_0_character_lcd_0_avalon_lcd_slave_write),                               //                                                         .write
		.character_lcd_0_avalon_lcd_slave_read                                (mm_interconnect_0_character_lcd_0_avalon_lcd_slave_read),                                //                                                         .read
		.character_lcd_0_avalon_lcd_slave_readdata                            (mm_interconnect_0_character_lcd_0_avalon_lcd_slave_readdata),                            //                                                         .readdata
		.character_lcd_0_avalon_lcd_slave_writedata                           (mm_interconnect_0_character_lcd_0_avalon_lcd_slave_writedata),                           //                                                         .writedata
		.character_lcd_0_avalon_lcd_slave_waitrequest                         (mm_interconnect_0_character_lcd_0_avalon_lcd_slave_waitrequest),                         //                                                         .waitrequest
		.character_lcd_0_avalon_lcd_slave_chipselect                          (mm_interconnect_0_character_lcd_0_avalon_lcd_slave_chipselect),                          //                                                         .chipselect
		.HEX_0_s1_address                                                     (mm_interconnect_0_hex_0_s1_address),                                                     //                                                 HEX_0_s1.address
		.HEX_0_s1_write                                                       (mm_interconnect_0_hex_0_s1_write),                                                       //                                                         .write
		.HEX_0_s1_readdata                                                    (mm_interconnect_0_hex_0_s1_readdata),                                                    //                                                         .readdata
		.HEX_0_s1_writedata                                                   (mm_interconnect_0_hex_0_s1_writedata),                                                   //                                                         .writedata
		.HEX_0_s1_chipselect                                                  (mm_interconnect_0_hex_0_s1_chipselect),                                                  //                                                         .chipselect
		.HEX_1_s1_address                                                     (mm_interconnect_0_hex_1_s1_address),                                                     //                                                 HEX_1_s1.address
		.HEX_1_s1_write                                                       (mm_interconnect_0_hex_1_s1_write),                                                       //                                                         .write
		.HEX_1_s1_readdata                                                    (mm_interconnect_0_hex_1_s1_readdata),                                                    //                                                         .readdata
		.HEX_1_s1_writedata                                                   (mm_interconnect_0_hex_1_s1_writedata),                                                   //                                                         .writedata
		.HEX_1_s1_chipselect                                                  (mm_interconnect_0_hex_1_s1_chipselect),                                                  //                                                         .chipselect
		.HEX_2_s1_address                                                     (mm_interconnect_0_hex_2_s1_address),                                                     //                                                 HEX_2_s1.address
		.HEX_2_s1_write                                                       (mm_interconnect_0_hex_2_s1_write),                                                       //                                                         .write
		.HEX_2_s1_readdata                                                    (mm_interconnect_0_hex_2_s1_readdata),                                                    //                                                         .readdata
		.HEX_2_s1_writedata                                                   (mm_interconnect_0_hex_2_s1_writedata),                                                   //                                                         .writedata
		.HEX_2_s1_chipselect                                                  (mm_interconnect_0_hex_2_s1_chipselect),                                                  //                                                         .chipselect
		.HEX_3_s1_address                                                     (mm_interconnect_0_hex_3_s1_address),                                                     //                                                 HEX_3_s1.address
		.HEX_3_s1_write                                                       (mm_interconnect_0_hex_3_s1_write),                                                       //                                                         .write
		.HEX_3_s1_readdata                                                    (mm_interconnect_0_hex_3_s1_readdata),                                                    //                                                         .readdata
		.HEX_3_s1_writedata                                                   (mm_interconnect_0_hex_3_s1_writedata),                                                   //                                                         .writedata
		.HEX_3_s1_chipselect                                                  (mm_interconnect_0_hex_3_s1_chipselect),                                                  //                                                         .chipselect
		.HEX_4_s1_address                                                     (mm_interconnect_0_hex_4_s1_address),                                                     //                                                 HEX_4_s1.address
		.HEX_4_s1_write                                                       (mm_interconnect_0_hex_4_s1_write),                                                       //                                                         .write
		.HEX_4_s1_readdata                                                    (mm_interconnect_0_hex_4_s1_readdata),                                                    //                                                         .readdata
		.HEX_4_s1_writedata                                                   (mm_interconnect_0_hex_4_s1_writedata),                                                   //                                                         .writedata
		.HEX_4_s1_chipselect                                                  (mm_interconnect_0_hex_4_s1_chipselect),                                                  //                                                         .chipselect
		.HEX_5_s1_address                                                     (mm_interconnect_0_hex_5_s1_address),                                                     //                                                 HEX_5_s1.address
		.HEX_5_s1_write                                                       (mm_interconnect_0_hex_5_s1_write),                                                       //                                                         .write
		.HEX_5_s1_readdata                                                    (mm_interconnect_0_hex_5_s1_readdata),                                                    //                                                         .readdata
		.HEX_5_s1_writedata                                                   (mm_interconnect_0_hex_5_s1_writedata),                                                   //                                                         .writedata
		.HEX_5_s1_chipselect                                                  (mm_interconnect_0_hex_5_s1_chipselect),                                                  //                                                         .chipselect
		.HEX_6_s1_address                                                     (mm_interconnect_0_hex_6_s1_address),                                                     //                                                 HEX_6_s1.address
		.HEX_6_s1_write                                                       (mm_interconnect_0_hex_6_s1_write),                                                       //                                                         .write
		.HEX_6_s1_readdata                                                    (mm_interconnect_0_hex_6_s1_readdata),                                                    //                                                         .readdata
		.HEX_6_s1_writedata                                                   (mm_interconnect_0_hex_6_s1_writedata),                                                   //                                                         .writedata
		.HEX_6_s1_chipselect                                                  (mm_interconnect_0_hex_6_s1_chipselect),                                                  //                                                         .chipselect
		.HEX_7_s1_address                                                     (mm_interconnect_0_hex_7_s1_address),                                                     //                                                 HEX_7_s1.address
		.HEX_7_s1_write                                                       (mm_interconnect_0_hex_7_s1_write),                                                       //                                                         .write
		.HEX_7_s1_readdata                                                    (mm_interconnect_0_hex_7_s1_readdata),                                                    //                                                         .readdata
		.HEX_7_s1_writedata                                                   (mm_interconnect_0_hex_7_s1_writedata),                                                   //                                                         .writedata
		.HEX_7_s1_chipselect                                                  (mm_interconnect_0_hex_7_s1_chipselect),                                                  //                                                         .chipselect
		.High_Res_Timer_s1_address                                            (mm_interconnect_0_high_res_timer_s1_address),                                            //                                        High_Res_Timer_s1.address
		.High_Res_Timer_s1_write                                              (mm_interconnect_0_high_res_timer_s1_write),                                              //                                                         .write
		.High_Res_Timer_s1_readdata                                           (mm_interconnect_0_high_res_timer_s1_readdata),                                           //                                                         .readdata
		.High_Res_Timer_s1_writedata                                          (mm_interconnect_0_high_res_timer_s1_writedata),                                          //                                                         .writedata
		.High_Res_Timer_s1_chipselect                                         (mm_interconnect_0_high_res_timer_s1_chipselect),                                         //                                                         .chipselect
		.jtag_uart_0_avalon_jtag_slave_address                                (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),                                //                            jtag_uart_0_avalon_jtag_slave.address
		.jtag_uart_0_avalon_jtag_slave_write                                  (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),                                  //                                                         .write
		.jtag_uart_0_avalon_jtag_slave_read                                   (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),                                   //                                                         .read
		.jtag_uart_0_avalon_jtag_slave_readdata                               (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),                               //                                                         .readdata
		.jtag_uart_0_avalon_jtag_slave_writedata                              (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),                              //                                                         .writedata
		.jtag_uart_0_avalon_jtag_slave_waitrequest                            (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest),                            //                                                         .waitrequest
		.jtag_uart_0_avalon_jtag_slave_chipselect                             (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),                             //                                                         .chipselect
		.KEY_0_s1_address                                                     (mm_interconnect_0_key_0_s1_address),                                                     //                                                 KEY_0_s1.address
		.KEY_0_s1_write                                                       (mm_interconnect_0_key_0_s1_write),                                                       //                                                         .write
		.KEY_0_s1_readdata                                                    (mm_interconnect_0_key_0_s1_readdata),                                                    //                                                         .readdata
		.KEY_0_s1_writedata                                                   (mm_interconnect_0_key_0_s1_writedata),                                                   //                                                         .writedata
		.KEY_0_s1_chipselect                                                  (mm_interconnect_0_key_0_s1_chipselect),                                                  //                                                         .chipselect
		.LEDG_s1_address                                                      (mm_interconnect_0_ledg_s1_address),                                                      //                                                  LEDG_s1.address
		.LEDG_s1_write                                                        (mm_interconnect_0_ledg_s1_write),                                                        //                                                         .write
		.LEDG_s1_readdata                                                     (mm_interconnect_0_ledg_s1_readdata),                                                     //                                                         .readdata
		.LEDG_s1_writedata                                                    (mm_interconnect_0_ledg_s1_writedata),                                                    //                                                         .writedata
		.LEDG_s1_chipselect                                                   (mm_interconnect_0_ledg_s1_chipselect),                                                   //                                                         .chipselect
		.LEDs_s1_address                                                      (mm_interconnect_0_leds_s1_address),                                                      //                                                  LEDs_s1.address
		.LEDs_s1_write                                                        (mm_interconnect_0_leds_s1_write),                                                        //                                                         .write
		.LEDs_s1_readdata                                                     (mm_interconnect_0_leds_s1_readdata),                                                     //                                                         .readdata
		.LEDs_s1_writedata                                                    (mm_interconnect_0_leds_s1_writedata),                                                    //                                                         .writedata
		.LEDs_s1_chipselect                                                   (mm_interconnect_0_leds_s1_chipselect),                                                   //                                                         .chipselect
		.myCPU_debug_mem_slave_address                                        (mm_interconnect_0_mycpu_debug_mem_slave_address),                                        //                                    myCPU_debug_mem_slave.address
		.myCPU_debug_mem_slave_write                                          (mm_interconnect_0_mycpu_debug_mem_slave_write),                                          //                                                         .write
		.myCPU_debug_mem_slave_read                                           (mm_interconnect_0_mycpu_debug_mem_slave_read),                                           //                                                         .read
		.myCPU_debug_mem_slave_readdata                                       (mm_interconnect_0_mycpu_debug_mem_slave_readdata),                                       //                                                         .readdata
		.myCPU_debug_mem_slave_writedata                                      (mm_interconnect_0_mycpu_debug_mem_slave_writedata),                                      //                                                         .writedata
		.myCPU_debug_mem_slave_byteenable                                     (mm_interconnect_0_mycpu_debug_mem_slave_byteenable),                                     //                                                         .byteenable
		.myCPU_debug_mem_slave_waitrequest                                    (mm_interconnect_0_mycpu_debug_mem_slave_waitrequest),                                    //                                                         .waitrequest
		.myCPU_debug_mem_slave_debugaccess                                    (mm_interconnect_0_mycpu_debug_mem_slave_debugaccess),                                    //                                                         .debugaccess
		.SDRAM_s1_address                                                     (mm_interconnect_0_sdram_s1_address),                                                     //                                                 SDRAM_s1.address
		.SDRAM_s1_write                                                       (mm_interconnect_0_sdram_s1_write),                                                       //                                                         .write
		.SDRAM_s1_read                                                        (mm_interconnect_0_sdram_s1_read),                                                        //                                                         .read
		.SDRAM_s1_readdata                                                    (mm_interconnect_0_sdram_s1_readdata),                                                    //                                                         .readdata
		.SDRAM_s1_writedata                                                   (mm_interconnect_0_sdram_s1_writedata),                                                   //                                                         .writedata
		.SDRAM_s1_byteenable                                                  (mm_interconnect_0_sdram_s1_byteenable),                                                  //                                                         .byteenable
		.SDRAM_s1_readdatavalid                                               (mm_interconnect_0_sdram_s1_readdatavalid),                                               //                                                         .readdatavalid
		.SDRAM_s1_waitrequest                                                 (mm_interconnect_0_sdram_s1_waitrequest),                                                 //                                                         .waitrequest
		.SDRAM_s1_chipselect                                                  (mm_interconnect_0_sdram_s1_chipselect),                                                  //                                                         .chipselect
		.Switches_s1_address                                                  (mm_interconnect_0_switches_s1_address),                                                  //                                              Switches_s1.address
		.Switches_s1_write                                                    (mm_interconnect_0_switches_s1_write),                                                    //                                                         .write
		.Switches_s1_readdata                                                 (mm_interconnect_0_switches_s1_readdata),                                                 //                                                         .readdata
		.Switches_s1_writedata                                                (mm_interconnect_0_switches_s1_writedata),                                                //                                                         .writedata
		.Switches_s1_chipselect                                               (mm_interconnect_0_switches_s1_chipselect),                                               //                                                         .chipselect
		.sysID_control_slave_address                                          (mm_interconnect_0_sysid_control_slave_address),                                          //                                      sysID_control_slave.address
		.sysID_control_slave_readdata                                         (mm_interconnect_0_sysid_control_slave_readdata),                                         //                                                         .readdata
		.System_Clock_Timer_s1_address                                        (mm_interconnect_0_system_clock_timer_s1_address),                                        //                                    System_Clock_Timer_s1.address
		.System_Clock_Timer_s1_write                                          (mm_interconnect_0_system_clock_timer_s1_write),                                          //                                                         .write
		.System_Clock_Timer_s1_readdata                                       (mm_interconnect_0_system_clock_timer_s1_readdata),                                       //                                                         .readdata
		.System_Clock_Timer_s1_writedata                                      (mm_interconnect_0_system_clock_timer_s1_writedata),                                      //                                                         .writedata
		.System_Clock_Timer_s1_chipselect                                     (mm_interconnect_0_system_clock_timer_s1_chipselect),                                     //                                                         .chipselect
		.TCM_s2_address                                                       (mm_interconnect_0_tcm_s2_address),                                                       //                                                   TCM_s2.address
		.TCM_s2_write                                                         (mm_interconnect_0_tcm_s2_write),                                                         //                                                         .write
		.TCM_s2_readdata                                                      (mm_interconnect_0_tcm_s2_readdata),                                                      //                                                         .readdata
		.TCM_s2_writedata                                                     (mm_interconnect_0_tcm_s2_writedata),                                                     //                                                         .writedata
		.TCM_s2_byteenable                                                    (mm_interconnect_0_tcm_s2_byteenable),                                                    //                                                         .byteenable
		.TCM_s2_chipselect                                                    (mm_interconnect_0_tcm_s2_chipselect),                                                    //                                                         .chipselect
		.TCM_s2_clken                                                         (mm_interconnect_0_tcm_s2_clken)                                                          //                                                         .clken
	);

	niosSys_mm_interconnect_1 mm_interconnect_1 (
		.MAIN_CLK_sys_clk_clk                                (main_clk_sys_clk_clk),                                //                           MAIN_CLK_sys_clk.clk
		.myCPU_reset_reset_bridge_in_reset_reset             (rst_controller_reset_out_reset),                      //          myCPU_reset_reset_bridge_in_reset.reset
		.myCPU_tightly_coupled_instruction_master_0_address  (mycpu_tightly_coupled_instruction_master_0_address),  // myCPU_tightly_coupled_instruction_master_0.address
		.myCPU_tightly_coupled_instruction_master_0_read     (mycpu_tightly_coupled_instruction_master_0_read),     //                                           .read
		.myCPU_tightly_coupled_instruction_master_0_readdata (mycpu_tightly_coupled_instruction_master_0_readdata), //                                           .readdata
		.myCPU_tightly_coupled_instruction_master_0_clken    (mycpu_tightly_coupled_instruction_master_0_clken),    //                                           .clken
		.TCM_s1_address                                      (mm_interconnect_1_tcm_s1_address),                    //                                     TCM_s1.address
		.TCM_s1_write                                        (mm_interconnect_1_tcm_s1_write),                      //                                           .write
		.TCM_s1_readdata                                     (mm_interconnect_1_tcm_s1_readdata),                   //                                           .readdata
		.TCM_s1_writedata                                    (mm_interconnect_1_tcm_s1_writedata),                  //                                           .writedata
		.TCM_s1_byteenable                                   (mm_interconnect_1_tcm_s1_byteenable),                 //                                           .byteenable
		.TCM_s1_chipselect                                   (mm_interconnect_1_tcm_s1_chipselect),                 //                                           .chipselect
		.TCM_s1_clken                                        (mm_interconnect_1_tcm_s1_clken)                       //                                           .clken
	);

	niosSys_irq_mapper irq_mapper (
		.clk           (main_clk_sys_clk_clk),           //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),       // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),       // receiver3.irq
		.receiver4_irq (irq_mapper_receiver4_irq),       // receiver4.irq
		.sender_irq    (mycpu_irq_irq)                   //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (mycpu_debug_reset_request_reset),    // reset_in0.reset
		.reset_in1      (main_clk_reset_source_reset),        // reset_in1.reset
		.clk            (main_clk_sys_clk_clk),               //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
